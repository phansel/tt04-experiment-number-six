module memory_chars(
input wire [9:0] addr,
output reg [15:0] dout //,
// input rst,
// input clk
);

//always @(posedge clk, posedge rst) begin
always @(addr) begin
    //if (rst)
    //    dout <= 16'b0010000000100000;
    case(addr) 
        10'b0000000000: dout <= 16'b0011000100110001;
        10'b0000000001: dout <= 16'b0010111100100000;
        10'b0000000010: dout <= 16'b0111001100100000;
        10'b0000000100: dout <= 16'b0010000000100000;
        10'b0000000101: dout <= 16'b0011000101110100;
        10'b0000000110: dout <= 16'b0010111100100000;
        10'b0000000111: dout <= 16'b0111001100100000;
        10'b0000001000: dout <= 16'b0101111000100000;
        10'b0000001001: dout <= 16'b0011001000100000;
        10'b0000001011: dout <= 16'b0010000000100000;
        10'b0000001100: dout <= 16'b0011000101110100;
        10'b0000001101: dout <= 16'b0010111101011110;
        10'b0000001110: dout <= 16'b0111001101111011;
        10'b0000001111: dout <= 16'b0101111001101110;
        10'b0000010000: dout <= 16'b0110111000101101;
        10'b0000010001: dout <= 16'b0010000000110001;
        10'b0000010010: dout <= 16'b0010000001111101;
        10'b0000010011: dout <= 16'b0010000000101111;
        10'b0000010100: dout <= 16'b0010000000101000;
        10'b0000010101: dout <= 16'b0010000001101110;
        10'b0000010110: dout <= 16'b0010000000101101;
        10'b0000010111: dout <= 16'b0010000000110001;
        10'b0000011000: dout <= 16'b0010000000101001;
        10'b0000011001: dout <= 16'b0010000000100001;
        10'b0000011011: dout <= 16'b0010000000100000;
        10'b0000011100: dout <= 16'b0011000100110001;
        10'b0000011101: dout <= 16'b0010111100101111;
        10'b0000011110: dout <= 16'b0101110001011100;
        10'b0000011111: dout <= 16'b0111001101110011;
        10'b0000100000: dout <= 16'b0111000101110001;
        10'b0000100001: dout <= 16'b0111001001110010;
        10'b0000100010: dout <= 16'b0111010001110100;
        10'b0000100011: dout <= 16'b0111101101111011;
        10'b0000100100: dout <= 16'b0111001101011100;
        10'b0000100101: dout <= 16'b0111110101110000;
        10'b0000100110: dout <= 16'b0010000001101001;
        10'b0000100111: dout <= 16'b0010000000100000;
        10'b0000101000: dout <= 16'b0010000001110100;
        10'b0000101001: dout <= 16'b0010000001111101;
        10'b0000101011: dout <= 16'b0010000000100000;
        10'b0000101100: dout <= 16'b0011000100110010;
        10'b0000101101: dout <= 16'b0010111101011100;
        10'b0000101110: dout <= 16'b0111001101110011;
        10'b0000101111: dout <= 16'b0101111001110001;
        10'b0000110000: dout <= 16'b0111101101110010;
        10'b0000110001: dout <= 16'b0011001101110100;
        10'b0000110010: dout <= 16'b0010111101111011;
        10'b0000110011: dout <= 16'b0011001001110100;
        10'b0000110100: dout <= 16'b0111110100101111;
        10'b0000110101: dout <= 16'b0010000001011100;
        10'b0000110110: dout <= 16'b0010000001110000;
        10'b0000110111: dout <= 16'b0010000001101001;
        10'b0000111000: dout <= 16'b0010000001111101;
        10'b0000111010: dout <= 16'b0010000000100000;
        10'b0000111011: dout <= 16'b0011000101110100;
        10'b0000111100: dout <= 16'b0010111101011110;
        10'b0000111101: dout <= 16'b0111001101111011;
        10'b0000111110: dout <= 16'b0101111001100001;
        10'b0000111111: dout <= 16'b0110000100101101;
        10'b0001000000: dout <= 16'b0010000000110001;
        10'b0001000001: dout <= 16'b0010000001111101;
        10'b0001000010: dout <= 16'b0010000000101111;
        10'b0001000011: dout <= 16'b0010000001011100;
        10'b0001000100: dout <= 16'b0010000001000111;
        10'b0001000101: dout <= 16'b0010000001100001;
        10'b0001000110: dout <= 16'b0010000001101101;
        10'b0001000111: dout <= 16'b0010000001101101;
        10'b0001001000: dout <= 16'b0010000001100001;
        10'b0001001001: dout <= 16'b0010000000101000;
        10'b0001001010: dout <= 16'b0010000001100001;
        10'b0001001011: dout <= 16'b0010000000101001;
        10'b0001001101: dout <= 16'b0010000000100000;
        10'b0001001110: dout <= 16'b0011000101100101;
        10'b0001001111: dout <= 16'b0010111101011110;
        10'b0001010000: dout <= 16'b0010100001111011;
        10'b0001010001: dout <= 16'b0111001101100001;
        10'b0001010010: dout <= 16'b0010110101110100;
        10'b0001010011: dout <= 16'b0110000101111101;
        10'b0001010100: dout <= 16'b0010100100100000;
        10'b0001010110: dout <= 16'b0010000000100000;
        10'b0001010111: dout <= 16'b0011000101110100;
        10'b0001011000: dout <= 16'b0010111101100101;
        10'b0001011001: dout <= 16'b0010100001011110;
        10'b0001011010: dout <= 16'b0111001101111011;
        10'b0001011011: dout <= 16'b0010110101100001;
        10'b0001011100: dout <= 16'b0110000101110100;
        10'b0001011101: dout <= 16'b0010100101111101;
        10'b0001011110: dout <= 16'b0101111000100000;
        10'b0001011111: dout <= 16'b0011001000100000;
        10'b0001100001: dout <= 16'b0010000000100000;
        10'b0001100010: dout <= 16'b0011000101011100;
        10'b0001100011: dout <= 16'b0010111101100110;
        10'b0001100100: dout <= 16'b0010100001110010;
        10'b0001100101: dout <= 16'b0111001101100001;
        10'b0001100110: dout <= 16'b0010110101100011;
        10'b0001100111: dout <= 16'b0110000101111011;
        10'b0001101000: dout <= 16'b0010100100110001;
        10'b0001101001: dout <= 16'b0101111001111101;
        10'b0001101010: dout <= 16'b0110111001111011;
        10'b0001101011: dout <= 16'b0010000000101000;
        10'b0001101100: dout <= 16'b0010000001101110;
        10'b0001101101: dout <= 16'b0010000000101101;
        10'b0001101110: dout <= 16'b0010000000110001;
        10'b0001101111: dout <= 16'b0010000000101001;
        10'b0001110000: dout <= 16'b0010000000100001;
        10'b0001110001: dout <= 16'b0010000001111101;
        10'b0001110010: dout <= 16'b0010000001110100;
        10'b0001110011: dout <= 16'b0010000001011110;
        10'b0001110100: dout <= 16'b0010000001111011;
        10'b0001110101: dout <= 16'b0010000001101110;
        10'b0001110110: dout <= 16'b0010000000101101;
        10'b0001110111: dout <= 16'b0010000000110001;
        10'b0001111000: dout <= 16'b0010000001111101;
        10'b0001111001: dout <= 16'b0010000001100101;
        10'b0001111010: dout <= 16'b0010000001011110;
        10'b0001111011: dout <= 16'b0010000001111011;
        10'b0001111100: dout <= 16'b0010000001100001;
        10'b0001111101: dout <= 16'b0010000001110100;
        10'b0001111110: dout <= 16'b0010000001111101;
        10'b0010000000: dout <= 16'b0010000000100000;
        10'b0010000001: dout <= 16'b0011000101011100;
        10'b0010000010: dout <= 16'b0010111101100110;
        10'b0010000011: dout <= 16'b0010100001110010;
        10'b0010000100: dout <= 16'b0111001101100001;
        10'b0010000101: dout <= 16'b0010110101100011;
        10'b0010000110: dout <= 16'b0110000101111011;
        10'b0010000111: dout <= 16'b0010100100110001;
        10'b0010001000: dout <= 16'b0101111001111101;
        10'b0010001001: dout <= 16'b0110101101111011;
        10'b0010001010: dout <= 16'b0010000001011100;
        10'b0010001011: dout <= 16'b0010000001000111;
        10'b0010001100: dout <= 16'b0010000001100001;
        10'b0010001101: dout <= 16'b0010000001101101;
        10'b0010001110: dout <= 16'b0010000001101101;
        10'b0010001111: dout <= 16'b0010000001100001;
        10'b0010010000: dout <= 16'b0010000000101000;
        10'b0010010001: dout <= 16'b0010000001101011;
        10'b0010010010: dout <= 16'b0010000000101001;
        10'b0010010011: dout <= 16'b0010000001111101;
        10'b0010010100: dout <= 16'b0010000001110100;
        10'b0010010101: dout <= 16'b0010000001011110;
        10'b0010010110: dout <= 16'b0010000001111011;
        10'b0010010111: dout <= 16'b0010000001101011;
        10'b0010011000: dout <= 16'b0010000000101101;
        10'b0010011001: dout <= 16'b0010000000110001;
        10'b0010011010: dout <= 16'b0010000001111101;
        10'b0010011011: dout <= 16'b0010000001100101;
        10'b0010011100: dout <= 16'b0010000001011110;
        10'b0010011101: dout <= 16'b0010000001111011;
        10'b0010011110: dout <= 16'b0010000001100001;
        10'b0010011111: dout <= 16'b0010000001110100;
        10'b0010100000: dout <= 16'b0010000001111101;
        10'b0010100010: dout <= 16'b0010000000100000;
        10'b0010100011: dout <= 16'b0101110001011100;
        10'b0010100100: dout <= 16'b0110011001100110;
        10'b0010100101: dout <= 16'b0111001001110010;
        10'b0010100110: dout <= 16'b0110000101100001;
        10'b0010100111: dout <= 16'b0110001101100011;
        10'b0010101000: dout <= 16'b0111101101111011;
        10'b0010101001: dout <= 16'b0011000100110001;
        10'b0010101010: dout <= 16'b0111110101111101;
        10'b0010101011: dout <= 16'b0111101101111011;
        10'b0010101100: dout <= 16'b0010100001100001;
        10'b0010101101: dout <= 16'b0111001100101101;
        10'b0010101110: dout <= 16'b0010110101100010;
        10'b0010101111: dout <= 16'b0110000101111101;
        10'b0010110000: dout <= 16'b0010100100101000;
        10'b0010110001: dout <= 16'b0010100001100101;
        10'b0010110010: dout <= 16'b0111001101011110;
        10'b0010110011: dout <= 16'b0010110101111011;
        10'b0010110100: dout <= 16'b0110001001100001;
        10'b0010110101: dout <= 16'b0010100101110100;
        10'b0010110110: dout <= 16'b0111110101111101;
        10'b0010110111: dout <= 16'b0010000000101101;
        10'b0010111000: dout <= 16'b0010000001100101;
        10'b0010111001: dout <= 16'b0010000001011110;
        10'b0010111010: dout <= 16'b0010000001111011;
        10'b0010111011: dout <= 16'b0010000001100010;
        10'b0010111100: dout <= 16'b0010000001110100;
        10'b0010111101: dout <= 16'b0010000001111101;
        10'b0010111110: dout <= 16'b0010000000101001;
        10'b0011000000: dout <= 16'b0010000000100000;
        10'b0011000001: dout <= 16'b0101110001011100;
        10'b0011000010: dout <= 16'b0110011001100110;
        10'b0011000011: dout <= 16'b0111001001110010;
        10'b0011000100: dout <= 16'b0110000101100001;
        10'b0011000101: dout <= 16'b0110001101100011;
        10'b0011000110: dout <= 16'b0111101101111011;
        10'b0011000111: dout <= 16'b0111001100110001;
        10'b0011001000: dout <= 16'b0111110101111101;
        10'b0011001001: dout <= 16'b0111101101111011;
        10'b0011001010: dout <= 16'b0010100001100001;
        10'b0011001011: dout <= 16'b0111001100101101;
        10'b0011001100: dout <= 16'b0010110101100010;
        10'b0011001101: dout <= 16'b0110000101111101;
        10'b0011001110: dout <= 16'b0010100100101000;
        10'b0011001111: dout <= 16'b0010100001100001;
        10'b0011010000: dout <= 16'b0111001101100101;
        10'b0011010001: dout <= 16'b0010110101011110;
        10'b0011010010: dout <= 16'b0110001001111011;
        10'b0011010011: dout <= 16'b0010100101100001;
        10'b0011010100: dout <= 16'b0111110101110100;
        10'b0011010101: dout <= 16'b0010000001111101;
        10'b0011010110: dout <= 16'b0010000000101101;
        10'b0011010111: dout <= 16'b0010000001100010;
        10'b0011011000: dout <= 16'b0010000001100101;
        10'b0011011001: dout <= 16'b0010000001011110;
        10'b0011011010: dout <= 16'b0010000001111011;
        10'b0011011011: dout <= 16'b0010000001100010;
        10'b0011011100: dout <= 16'b0010000001110100;
        10'b0011011101: dout <= 16'b0010000001111101;
        10'b0011011110: dout <= 16'b0010000000101001;
        10'b0011100000: dout <= 16'b0010000000100000;
        10'b0011100001: dout <= 16'b0101110001011100;
        10'b0011100010: dout <= 16'b0110011001100110;
        10'b0011100011: dout <= 16'b0111001001110010;
        10'b0011100100: dout <= 16'b0110000101100001;
        10'b0011100101: dout <= 16'b0110001101100011;
        10'b0011100110: dout <= 16'b0111101101111011;
        10'b0011100111: dout <= 16'b0011000100110001;
        10'b0011101000: dout <= 16'b0111110101111101;
        10'b0011101001: dout <= 16'b0111101101111011;
        10'b0011101010: dout <= 16'b0111001101011100;
        10'b0011101011: dout <= 16'b0101111001101111;
        10'b0011101100: dout <= 16'b0011001001101101;
        10'b0011101101: dout <= 16'b0010101101100101;
        10'b0011101110: dout <= 16'b0101110001100111;
        10'b0011101111: dout <= 16'b0110111101100001;
        10'b0011110000: dout <= 16'b0110110101111101;
        10'b0011110001: dout <= 16'b0110010101011100;
        10'b0011110010: dout <= 16'b0110011101110011;
        10'b0011110011: dout <= 16'b0110000101101001;
        10'b0011110100: dout <= 16'b0101111001101110;
        10'b0011110101: dout <= 16'b0011001000100000;
        10'b0011110110: dout <= 16'b0111110101011100;
        10'b0011110111: dout <= 16'b0010000001101111;
        10'b0011111000: dout <= 16'b0010000001101101;
        10'b0011111001: dout <= 16'b0010000001100101;
        10'b0011111010: dout <= 16'b0010000001100111;
        10'b0011111011: dout <= 16'b0010000001100001;
        10'b0011111100: dout <= 16'b0010000000100000;
        10'b0011111101: dout <= 16'b0010000001110100;
        10'b0011111111: dout <= 16'b0010000000100000;
        10'b0100000000: dout <= 16'b0101110001011100;
        10'b0100000001: dout <= 16'b0110011001100011;
        10'b0100000010: dout <= 16'b0111001001101111;
        10'b0100000011: dout <= 16'b0110000101110011;
        10'b0100000100: dout <= 16'b0110001100100000;
        10'b0100000101: dout <= 16'b0111101101011100;
        10'b0100000110: dout <= 16'b0111001101101111;
        10'b0100000111: dout <= 16'b0111110101101101;
        10'b0100001000: dout <= 16'b0111101101100101;
        10'b0100001001: dout <= 16'b0111001101100111;
        10'b0100001010: dout <= 16'b0101111001100001;
        10'b0100001011: dout <= 16'b0011001000100000;
        10'b0100001100: dout <= 16'b0010101100100000;
        10'b0100001101: dout <= 16'b0101110000100000;
        10'b0100001110: dout <= 16'b0110111100100000;
        10'b0100001111: dout <= 16'b0110110100100000;
        10'b0100010000: dout <= 16'b0110010100100000;
        10'b0100010001: dout <= 16'b0110011100100000;
        10'b0100010010: dout <= 16'b0110000100100000;
        10'b0100010011: dout <= 16'b0101111000100000;
        10'b0100010100: dout <= 16'b0011001000100000;
        10'b0100010101: dout <= 16'b0111110100100000;
        10'b0100010111: dout <= 16'b0010000000100000;
        10'b0100011000: dout <= 16'b0101110001011100;
        10'b0100011001: dout <= 16'b0110011001100110;
        10'b0100011010: dout <= 16'b0111001001110010;
        10'b0100011011: dout <= 16'b0110000101100001;
        10'b0100011100: dout <= 16'b0110001101100011;
        10'b0100011101: dout <= 16'b0111101101111011;
        10'b0100011110: dout <= 16'b0011000100110001;
        10'b0100011111: dout <= 16'b0111110101111101;
        10'b0100100000: dout <= 16'b0111101101111011;
        10'b0100100001: dout <= 16'b0111001101100001;
        10'b0100100010: dout <= 16'b0101111001111101;
        10'b0100100011: dout <= 16'b0011001001011100;
        10'b0100100100: dout <= 16'b0010110101110011;
        10'b0100100101: dout <= 16'b0110000101101001;
        10'b0100100110: dout <= 16'b0101111001101110;
        10'b0100100111: dout <= 16'b0011001001101000;
        10'b0100101000: dout <= 16'b0111110100100000;
        10'b0100101001: dout <= 16'b0010000001100001;
        10'b0100101010: dout <= 16'b0010000001110100;
        10'b0100101100: dout <= 16'b0010000000100000;
        10'b0100101101: dout <= 16'b0101110001011100;
        10'b0100101110: dout <= 16'b0110011001100011;
        10'b0100101111: dout <= 16'b0111001001101111;
        10'b0100110000: dout <= 16'b0110000101110011;
        10'b0100110001: dout <= 16'b0110001101101000;
        10'b0100110010: dout <= 16'b0111101100100000;
        10'b0100110011: dout <= 16'b0111001101100001;
        10'b0100110100: dout <= 16'b0111110101110100;
        10'b0100110101: dout <= 16'b0111101100100000;
        10'b0100110110: dout <= 16'b0111001100100000;
        10'b0100110111: dout <= 16'b0101111000100000;
        10'b0100111000: dout <= 16'b0011001000100000;
        10'b0100111001: dout <= 16'b0010110100100000;
        10'b0100111010: dout <= 16'b0110000100100000;
        10'b0100111011: dout <= 16'b0101111000100000;
        10'b0100111100: dout <= 16'b0011001000100000;
        10'b0100111101: dout <= 16'b0111110100100000;
        10'b0100111111: dout <= 16'b0010000000100000;
        10'b0101000000: dout <= 16'b0101110001011100;
        10'b0101000001: dout <= 16'b0110011001100110;
        10'b0101000010: dout <= 16'b0111001001110010;
        10'b0101000011: dout <= 16'b0110000101100001;
        10'b0101000100: dout <= 16'b0110001101100011;
        10'b0101000101: dout <= 16'b0111101101111011;
        10'b0101000110: dout <= 16'b0011000100110001;
        10'b0101000111: dout <= 16'b0111110101111101;
        10'b0101001000: dout <= 16'b0111101101111011;
        10'b0101001001: dout <= 16'b0010100001011100;
        10'b0101001010: dout <= 16'b0111001101101111;
        10'b0101001011: dout <= 16'b0010110101101101;
        10'b0101001100: dout <= 16'b0110000101100101;
        10'b0101001101: dout <= 16'b0010100101100111;
        10'b0101001110: dout <= 16'b0101111001100001;
        10'b0101001111: dout <= 16'b0011001001111101;
        10'b0101010000: dout <= 16'b0010101100100000;
        10'b0101010001: dout <= 16'b0101110001100101;
        10'b0101010010: dout <= 16'b0110111101011110;
        10'b0101010011: dout <= 16'b0110110101111011;
        10'b0101010100: dout <= 16'b0110010101100001;
        10'b0101010101: dout <= 16'b0110011101110100;
        10'b0101010110: dout <= 16'b0110000101111101;
        10'b0101010111: dout <= 16'b0101111001011100;
        10'b0101011000: dout <= 16'b0011001001110011;
        10'b0101011001: dout <= 16'b0111110101101001;
        10'b0101011010: dout <= 16'b0010000001101110;
        10'b0101011011: dout <= 16'b0010000001101000;
        10'b0101011100: dout <= 16'b0010000000100000;
        10'b0101011101: dout <= 16'b0010000001011100;
        10'b0101011110: dout <= 16'b0010000001101111;
        10'b0101011111: dout <= 16'b0010000001101101;
        10'b0101100000: dout <= 16'b0010000001100101;
        10'b0101100001: dout <= 16'b0010000001100111;
        10'b0101100010: dout <= 16'b0010000001100001;
        10'b0101100011: dout <= 16'b0010000000100000;
        10'b0101100100: dout <= 16'b0010000001110100;
        10'b0101100110: dout <= 16'b0010000000100000;
        10'b0101100111: dout <= 16'b0101110001100101;
        10'b0101101000: dout <= 16'b0110011001011110;
        10'b0101101001: dout <= 16'b0111001001111011;
        10'b0101101010: dout <= 16'b0110000101100001;
        10'b0101101011: dout <= 16'b0110001101110100;
        10'b0101101100: dout <= 16'b0111101101111101;
        10'b0101101101: dout <= 16'b0111001101011100;
        10'b0101101110: dout <= 16'b0010110101100011;
        10'b0101101111: dout <= 16'b0110000101101111;
        10'b0101110000: dout <= 16'b0111110101110011;
        10'b0101110001: dout <= 16'b0111101100100000;
        10'b0101110010: dout <= 16'b0010100001011100;
        10'b0101110011: dout <= 16'b0111001101101111;
        10'b0101110100: dout <= 16'b0010110101101101;
        10'b0101110101: dout <= 16'b0110000101100101;
        10'b0101110110: dout <= 16'b0010100101100111;
        10'b0101110111: dout <= 16'b0101111001100001;
        10'b0101111000: dout <= 16'b0011001000100000;
        10'b0101111001: dout <= 16'b0010000001110100;
        10'b0101111010: dout <= 16'b0010101100100000;
        10'b0101111011: dout <= 16'b0010000000100000;
        10'b0101111100: dout <= 16'b0101110000100000;
        10'b0101111101: dout <= 16'b0110111100100000;
        10'b0101111110: dout <= 16'b0110110100100000;
        10'b0101111111: dout <= 16'b0110010100100000;
        10'b0110000000: dout <= 16'b0110011100100000;
        10'b0110000001: dout <= 16'b0110000100100000;
        10'b0110000010: dout <= 16'b0101111000100000;
        10'b0110000011: dout <= 16'b0011001000100000;
        10'b0110000100: dout <= 16'b0111110100100000;
        10'b0110000110: dout <= 16'b0010000000100000;
        10'b0110000111: dout <= 16'b0101110001011100;
        10'b0110001000: dout <= 16'b0110011001100110;
        10'b0110001001: dout <= 16'b0111001001110010;
        10'b0110001010: dout <= 16'b0110000101100001;
        10'b0110001011: dout <= 16'b0110001101100011;
        10'b0110001100: dout <= 16'b0111101101111011;
        10'b0110001101: dout <= 16'b0011000100110001;
        10'b0110001110: dout <= 16'b0111110101111101;
        10'b0110001111: dout <= 16'b0111101101111011;
        10'b0110010000: dout <= 16'b0111001101011100;
        10'b0110010001: dout <= 16'b0010100001101111;
        10'b0110010010: dout <= 16'b0111001101101101;
        10'b0110010011: dout <= 16'b0101111001100101;
        10'b0110010100: dout <= 16'b0111001101100111;
        10'b0110010101: dout <= 16'b0010101101100001;
        10'b0110010110: dout <= 16'b0101110001011110;
        10'b0110010111: dout <= 16'b0110111100110010;
        10'b0110011000: dout <= 16'b0110110101111101;
        10'b0110011001: dout <= 16'b0110010100101000;
        10'b0110011010: dout <= 16'b0110011100110001;
        10'b0110011011: dout <= 16'b0110000100101101;
        10'b0110011100: dout <= 16'b0101111001011100;
        10'b0110011101: dout <= 16'b0011001001100011;
        10'b0110011110: dout <= 16'b0111110101101111;
        10'b0110011111: dout <= 16'b0010000001110011;
        10'b0110100000: dout <= 16'b0010000000100000;
        10'b0110100001: dout <= 16'b0010000001011100;
        10'b0110100010: dout <= 16'b0010000001101111;
        10'b0110100011: dout <= 16'b0010000001101101;
        10'b0110100100: dout <= 16'b0010000001100101;
        10'b0110100101: dout <= 16'b0010000001100111;
        10'b0110100110: dout <= 16'b0010000001100001;
        10'b0110100111: dout <= 16'b0010000000100000;
        10'b0110101000: dout <= 16'b0010000001110100;
        10'b0110101001: dout <= 16'b0010000000101001;
        10'b0110101011: dout <= 16'b0010000000100000;
        10'b0110101100: dout <= 16'b0101110001011100;
        10'b0110101101: dout <= 16'b0110011001100110;
        10'b0110101110: dout <= 16'b0111001001110010;
        10'b0110101111: dout <= 16'b0110000101100001;
        10'b0110110000: dout <= 16'b0110001101100011;
        10'b0110110001: dout <= 16'b0111101101111011;
        10'b0110110010: dout <= 16'b0011000100110001;
        10'b0110110011: dout <= 16'b0111110101111101;
        10'b0110110100: dout <= 16'b0111101101111011;
        10'b0110110101: dout <= 16'b0111001101011100;
        10'b0110110110: dout <= 16'b0101111001101111;
        10'b0110110111: dout <= 16'b0011001001101101;
        10'b0110111000: dout <= 16'b0010100001100101;
        10'b0110111001: dout <= 16'b0111001101100111;
        10'b0110111010: dout <= 16'b0101111001100001;
        10'b0110111011: dout <= 16'b0011001001011110;
        10'b0110111100: dout <= 16'b0010101100110011;
        10'b0110111101: dout <= 16'b0101110001111101;
        10'b0110111110: dout <= 16'b0110111100101000;
        10'b0110111111: dout <= 16'b0110110101011100;
        10'b0111000000: dout <= 16'b0110010101101111;
        10'b0111000001: dout <= 16'b0110011101101101;
        10'b0111000010: dout <= 16'b0110000101100101;
        10'b0111000011: dout <= 16'b0101111001100111;
        10'b0111000100: dout <= 16'b0011001001100001;
        10'b0111000101: dout <= 16'b0010100100100000;
        10'b0111000110: dout <= 16'b0111110101110100;
        10'b0111000111: dout <= 16'b0010000000100000;
        10'b0111001000: dout <= 16'b0010000000101101;
        10'b0111001001: dout <= 16'b0010000000100000;
        10'b0111001010: dout <= 16'b0010000001011100;
        10'b0111001011: dout <= 16'b0010000001110011;
        10'b0111001100: dout <= 16'b0010000001101001;
        10'b0111001101: dout <= 16'b0010000001101110;
        10'b0111001110: dout <= 16'b0010000000100000;
        10'b0111001111: dout <= 16'b0010000001011100;
        10'b0111010000: dout <= 16'b0010000001101111;
        10'b0111010001: dout <= 16'b0010000001101101;
        10'b0111010010: dout <= 16'b0010000001100101;
        10'b0111010011: dout <= 16'b0010000001100111;
        10'b0111010100: dout <= 16'b0010000001100001;
        10'b0111010101: dout <= 16'b0010000000100000;
        10'b0111010110: dout <= 16'b0010000001110100;
        10'b0111010111: dout <= 16'b0010000000101001;
        10'b0111011001: dout <= 16'b0010000000100000;
        10'b0111011010: dout <= 16'b0101110001011100;
        10'b0111011011: dout <= 16'b0110011001100110;
        10'b0111011100: dout <= 16'b0111001001110010;
        10'b0111011101: dout <= 16'b0110000101100001;
        10'b0111011110: dout <= 16'b0110001101100011;
        10'b0111011111: dout <= 16'b0111101101111011;
        10'b0111100000: dout <= 16'b0011000100110001;
        10'b0111100001: dout <= 16'b0111110101111101;
        10'b0111100010: dout <= 16'b0111101101111011;
        10'b0111100011: dout <= 16'b0010100000110010;
        10'b0111100100: dout <= 16'b0111001101011100;
        10'b0111100101: dout <= 16'b0101111001101111;
        10'b0111100110: dout <= 16'b0011001001101101;
        10'b0111100111: dout <= 16'b0010101101100101;
        10'b0111101000: dout <= 16'b0101110001100111;
        10'b0111101001: dout <= 16'b0110111101100001;
        10'b0111101010: dout <= 16'b0110110101011110;
        10'b0111101011: dout <= 16'b0110010100110011;
        10'b0111101100: dout <= 16'b0110011101111101;
        10'b0111101101: dout <= 16'b0110000100101000;
        10'b0111101110: dout <= 16'b0101111001011100;
        10'b0111101111: dout <= 16'b0011001001110011;
        10'b0111110000: dout <= 16'b0010100101101001;
        10'b0111110001: dout <= 16'b0101111001101110;
        10'b0111110010: dout <= 16'b0011001000100000;
        10'b0111110011: dout <= 16'b0111110101011100;
        10'b0111110100: dout <= 16'b0010000001101111;
        10'b0111110101: dout <= 16'b0010000001101101;
        10'b0111110110: dout <= 16'b0010000001100101;
        10'b0111110111: dout <= 16'b0010000001100111;
        10'b0111111000: dout <= 16'b0010000001100001;
        10'b0111111001: dout <= 16'b0010000000100000;
        10'b0111111010: dout <= 16'b0010000001110100;
        10'b0111111011: dout <= 16'b0010000000100000;
        10'b0111111100: dout <= 16'b0010000000101101;
        10'b0111111101: dout <= 16'b0010000000100000;
        10'b0111111110: dout <= 16'b0010000001011100;
        10'b0111111111: dout <= 16'b0010000001101111;
        10'b1000000000: dout <= 16'b0010000001101101;
        10'b1000000001: dout <= 16'b0010000001100101;
        10'b1000000010: dout <= 16'b0010000001100111;
        10'b1000000011: dout <= 16'b0010000001100001;
        10'b1000000100: dout <= 16'b0010000000100000;
        10'b1000000101: dout <= 16'b0010000001110100;
        10'b1000000110: dout <= 16'b0010000000100000;
        10'b1000000111: dout <= 16'b0010000001011100;
        10'b1000001000: dout <= 16'b0010000001100011;
        10'b1000001001: dout <= 16'b0010000001101111;
        10'b1000001010: dout <= 16'b0010000001110011;
        10'b1000001011: dout <= 16'b0010000000100000;
        10'b1000001100: dout <= 16'b0010000001011100;
        10'b1000001101: dout <= 16'b0010000001101111;
        10'b1000001110: dout <= 16'b0010000001101101;
        10'b1000001111: dout <= 16'b0010000001100101;
        10'b1000010000: dout <= 16'b0010000001100111;
        10'b1000010001: dout <= 16'b0010000001100001;
        10'b1000010010: dout <= 16'b0010000000100000;
        10'b1000010011: dout <= 16'b0010000001110100;
        10'b1000010100: dout <= 16'b0010000000101001;
        10'b1000010110: dout <= 16'b0010000000100000;
        10'b1000010111: dout <= 16'b0101110001011100;
        10'b1000011000: dout <= 16'b0110011001100110;
        10'b1000011001: dout <= 16'b0111001001110010;
        10'b1000011010: dout <= 16'b0110000101100001;
        10'b1000011011: dout <= 16'b0110001101100011;
        10'b1000011100: dout <= 16'b0111101101111011;
        10'b1000011101: dout <= 16'b0111001100110001;
        10'b1000011110: dout <= 16'b0111110101111101;
        10'b1000011111: dout <= 16'b0111101101111011;
        10'b1000100000: dout <= 16'b0010100000110010;
        10'b1000100001: dout <= 16'b0111001101011100;
        10'b1000100010: dout <= 16'b0101111001101111;
        10'b1000100011: dout <= 16'b0011001001101101;
        10'b1000100100: dout <= 16'b0010101101100101;
        10'b1000100101: dout <= 16'b0101110001100111;
        10'b1000100110: dout <= 16'b0110111101100001;
        10'b1000100111: dout <= 16'b0110110101111101;
        10'b1000101000: dout <= 16'b0110010101011100;
        10'b1000101001: dout <= 16'b0110011101110011;
        10'b1000101010: dout <= 16'b0110000101101001;
        10'b1000101011: dout <= 16'b0101111001101110;
        10'b1000101100: dout <= 16'b0011001000100000;
        10'b1000101101: dout <= 16'b0010100101011100;
        10'b1000101110: dout <= 16'b0101111001101111;
        10'b1000101111: dout <= 16'b0011001001101101;
        10'b1000110000: dout <= 16'b0111110101100101;
        10'b1000110001: dout <= 16'b0010000001100111;
        10'b1000110010: dout <= 16'b0010000001100001;
        10'b1000110011: dout <= 16'b0010000000100000;
        10'b1000110100: dout <= 16'b0010000001110100;
        10'b1000110110: dout <= 16'b0010000000100000;
        10'b1000110111: dout <= 16'b0101110001011100;
        10'b1000111000: dout <= 16'b0110011001100110;
        10'b1000111001: dout <= 16'b0111001001110010;
        10'b1000111010: dout <= 16'b0110000101100001;
        10'b1000111011: dout <= 16'b0110001101100011;
        10'b1000111100: dout <= 16'b0111101101111011;
        10'b1000111101: dout <= 16'b0111001100110001;
        10'b1000111110: dout <= 16'b0101111001111101;
        10'b1000111111: dout <= 16'b0011001001111011;
        10'b1001000000: dout <= 16'b0111110100110010;
        10'b1001000001: dout <= 16'b0111101101011100;
        10'b1001000010: dout <= 16'b0010100001101111;
        10'b1001000011: dout <= 16'b0111001101101101;
        10'b1001000100: dout <= 16'b0101111001100101;
        10'b1001000101: dout <= 16'b0011001001100111;
        10'b1001000110: dout <= 16'b0010101101100001;
        10'b1001000111: dout <= 16'b0101110001111101;
        10'b1001001000: dout <= 16'b0110111100101000;
        10'b1001001001: dout <= 16'b0110110101011100;
        10'b1001001010: dout <= 16'b0110010101110011;
        10'b1001001011: dout <= 16'b0110011101101001;
        10'b1001001100: dout <= 16'b0110000101101110;
        10'b1001001101: dout <= 16'b0101111000100000;
        10'b1001001110: dout <= 16'b0011001001011100;
        10'b1001001111: dout <= 16'b0010100101101111;
        10'b1001010000: dout <= 16'b0101111001101101;
        10'b1001010001: dout <= 16'b0011001001100101;
        10'b1001010010: dout <= 16'b0111110101100111;
        10'b1001010011: dout <= 16'b0010000001100001;
        10'b1001010100: dout <= 16'b0010000000100000;
        10'b1001010101: dout <= 16'b0010000001110100;
        10'b1001010110: dout <= 16'b0010000000101011;
        10'b1001010111: dout <= 16'b0010000001011100;
        10'b1001011000: dout <= 16'b0010000001101111;
        10'b1001011001: dout <= 16'b0010000001101101;
        10'b1001011010: dout <= 16'b0010000001100101;
        10'b1001011011: dout <= 16'b0010000001100111;
        10'b1001011100: dout <= 16'b0010000001100001;
        10'b1001011101: dout <= 16'b0010000000100000;
        10'b1001011110: dout <= 16'b0010000001110100;
        10'b1001011111: dout <= 16'b0010000001011100;
        10'b1001100000: dout <= 16'b0010000001100011;
        10'b1001100001: dout <= 16'b0010000001101111;
        10'b1001100010: dout <= 16'b0010000001110011;
        10'b1001100011: dout <= 16'b0010000001011100;
        10'b1001100100: dout <= 16'b0010000001101111;
        10'b1001100101: dout <= 16'b0010000001101101;
        10'b1001100110: dout <= 16'b0010000001100101;
        10'b1001100111: dout <= 16'b0010000001100111;
        10'b1001101000: dout <= 16'b0010000001100001;
        10'b1001101001: dout <= 16'b0010000000100000;
        10'b1001101010: dout <= 16'b0010000001110100;
        10'b1001101011: dout <= 16'b0010000000101001;
        10'b1001101101: dout <= 16'b0010000000100000;
        10'b1001101110: dout <= 16'b0101110001011100;
        10'b1001101111: dout <= 16'b0110011001100110;
        10'b1001110000: dout <= 16'b0111001001110010;
        10'b1001110001: dout <= 16'b0110000101100001;
        10'b1001110010: dout <= 16'b0110001101100011;
        10'b1001110011: dout <= 16'b0111101101111011;
        10'b1001110100: dout <= 16'b0111001100110001;
        10'b1001110101: dout <= 16'b0111110101111101;
        10'b1001110110: dout <= 16'b0111101101111011;
        10'b1001110111: dout <= 16'b0010100001100010;
        10'b1001111000: dout <= 16'b0111001101011110;
        10'b1001111001: dout <= 16'b0101111000110010;
        10'b1001111010: dout <= 16'b0011001000101101;
        10'b1001111011: dout <= 16'b0010101101100001;
        10'b1001111100: dout <= 16'b0110000101011110;
        10'b1001111101: dout <= 16'b0101111000110010;
        10'b1001111110: dout <= 16'b0011001001111101;
        10'b1001111111: dout <= 16'b0010100100101000;
        10'b1010000000: dout <= 16'b0010100001011100;
        10'b1010000001: dout <= 16'b0111001101100011;
        10'b1010000010: dout <= 16'b0101111001101111;
        10'b1010000011: dout <= 16'b0011001001110011;
        10'b1010000100: dout <= 16'b0010101100100000;
        10'b1010000101: dout <= 16'b0110001001100001;
        10'b1010000110: dout <= 16'b0101111001110100;
        10'b1010000111: dout <= 16'b0011001000101101;
        10'b1010001000: dout <= 16'b0010100101011100;
        10'b1010001001: dout <= 16'b0111110101100011;
        10'b1010001010: dout <= 16'b0010000001101111;
        10'b1010001011: dout <= 16'b0010000001110011;
        10'b1010001100: dout <= 16'b0010000000100000;
        10'b1010001101: dout <= 16'b0010000001100010;
        10'b1010001110: dout <= 16'b0010000001110100;
        10'b1010001111: dout <= 16'b0010000000101001;
        10'b1010010001: dout <= 16'b0010000000100000;
        default: dout <= 16'b0010000000100000;
    endcase;
end

endmodule



module line_mapper(
//input wire clk,
//input wire rst,
input wire [7:0] line, 
output reg [19:0] addr);

//always @(posedge clk, posedge rst) begin
always @(line) begin
    // if (rst)
    //     addr <= 20'b000000011000000000;
    case(line)
    8'b00000000: addr <= 20'b00000000110000000000;
    8'b00000001: addr <= 20'b00000001010000000101;
    8'b00000010: addr <= 20'b00000011100000001100;
    8'b00000011: addr <= 20'b00000011100000011100;
    8'b00000100: addr <= 20'b00000011010000101100;
    8'b00000101: addr <= 20'b00000100010000111011;
    8'b00000110: addr <= 20'b00000001110001001110;
    8'b00000111: addr <= 20'b00000010010001010111;
    8'b00001000: addr <= 20'b00000111010001100010;
    8'b00001001: addr <= 20'b00001000000010000001;
    8'b00001010: addr <= 20'b00000111000010100011;
    8'b00001011: addr <= 20'b00000111100011000001;
    8'b00001100: addr <= 20'b00000111010011100001;
    8'b00001101: addr <= 20'b00000101100100000000;
    8'b00001110: addr <= 20'b00000100110100011000;
    8'b00001111: addr <= 20'b00000100010100101101;
    8'b00010000: addr <= 20'b00001001010101000000;
    8'b00010001: addr <= 20'b00000111100101100111;
    8'b00010010: addr <= 20'b00001000110110000111;
    8'b00010011: addr <= 20'b00001011000110101100;
    8'b00010100: addr <= 20'b00001110110111011010;
    8'b00010101: addr <= 20'b00000111101000010111;
    8'b00010110: addr <= 20'b00001101011000110111;
    8'b00010111: addr <= 20'b00001000101001101110;
    default: addr <= 20'b00000000110000000000;
    endcase;
end

endmodule



