module memory_chars(
input wire [7:0] addr, 
output reg [15:0] dout //,
// input rst,
// input clk
);

//always @(posedge clk, posedge rst) begin
always @(addr) begin
    //if (rst)
    //    dout <= 16'b0010000000100000;
    case(addr) 
        8'b00000000: dout <= 16'b0011000100110001;
        8'b00000001: dout <= 16'b0010111100100000;
        8'b00000010: dout <= 16'b0111001100100000;
        8'b00000100: dout <= 16'b0010000000100000;
        8'b00000101: dout <= 16'b0011000101110100;
        8'b00000110: dout <= 16'b0010111100100000;
        8'b00000111: dout <= 16'b0111001100100000;
        8'b00001000: dout <= 16'b0101111000100000;
        8'b00001001: dout <= 16'b0011001000100000;
        8'b00001011: dout <= 16'b0010000000100000;
        8'b00001100: dout <= 16'b0011000101110100;
        8'b00001101: dout <= 16'b0010111101011110;
        8'b00001110: dout <= 16'b0111001101111011;
        8'b00001111: dout <= 16'b0101111001101110;
        8'b00010000: dout <= 16'b0110111000101101;
        8'b00010001: dout <= 16'b0010000000110001;
        8'b00010010: dout <= 16'b0010000001111101;
        8'b00010011: dout <= 16'b0010000000101111;
        8'b00010100: dout <= 16'b0010000000101000;
        8'b00010101: dout <= 16'b0010000001101110;
        8'b00010110: dout <= 16'b0010000000101101;
        8'b00010111: dout <= 16'b0010000000110001;
        8'b00011000: dout <= 16'b0010000000101001;
        8'b00011001: dout <= 16'b0010000000100001;
        8'b00011011: dout <= 16'b0010000000100000;
        8'b00011100: dout <= 16'b0011000100110001;
        8'b00011101: dout <= 16'b0010111100101111;
        8'b00011110: dout <= 16'b0101110001011100;
        8'b00011111: dout <= 16'b0111001101110011;
        8'b00100000: dout <= 16'b0111000101110001;
        8'b00100001: dout <= 16'b0111001001110010;
        8'b00100010: dout <= 16'b0111010001110100;
        8'b00100011: dout <= 16'b0111101101111011;
        8'b00100100: dout <= 16'b0111001101011100;
        8'b00100101: dout <= 16'b0111110101110000;
        8'b00100110: dout <= 16'b0010000001101001;
        8'b00100111: dout <= 16'b0010000000100000;
        8'b00101000: dout <= 16'b0010000001110100;
        8'b00101001: dout <= 16'b0010000001111101;
        8'b00101011: dout <= 16'b0010000000100000;
        8'b00101100: dout <= 16'b0011000100110010;
        8'b00101101: dout <= 16'b0010111101011100;
        8'b00101110: dout <= 16'b0111001101110011;
        8'b00101111: dout <= 16'b0101111001110001;
        8'b00110000: dout <= 16'b0111101101110010;
        8'b00110001: dout <= 16'b0011001101110100;
        8'b00110010: dout <= 16'b0010111101111011;
        8'b00110011: dout <= 16'b0011001001110100;
        8'b00110100: dout <= 16'b0111110100101111;
        8'b00110101: dout <= 16'b0010000001011100;
        8'b00110110: dout <= 16'b0010000001110000;
        8'b00110111: dout <= 16'b0010000001101001;
        8'b00111000: dout <= 16'b0010000001111101;
        8'b00111010: dout <= 16'b0010000000100000;
        8'b00111011: dout <= 16'b0011000101110100;
        8'b00111100: dout <= 16'b0010111101011110;
        8'b00111101: dout <= 16'b0111001101111011;
        8'b00111110: dout <= 16'b0101111001100001;
        8'b00111111: dout <= 16'b0110000100101101;
        8'b01000000: dout <= 16'b0010000000110001;
        8'b01000001: dout <= 16'b0010000001111101;
        8'b01000010: dout <= 16'b0010000000101111;
        8'b01000011: dout <= 16'b0010000001011100;
        8'b01000100: dout <= 16'b0010000001000111;
        8'b01000101: dout <= 16'b0010000001100001;
        8'b01000110: dout <= 16'b0010000001101101;
        8'b01000111: dout <= 16'b0010000001101101;
        8'b01001000: dout <= 16'b0010000001100001;
        8'b01001001: dout <= 16'b0010000000101000;
        8'b01001010: dout <= 16'b0010000001100001;
        8'b01001011: dout <= 16'b0010000000101001;
        8'b01001101: dout <= 16'b0010000000100000;
        8'b01001110: dout <= 16'b0011000101100101;
        8'b01001111: dout <= 16'b0010111101011110;
        8'b01010000: dout <= 16'b0010100001111011;
        8'b01010001: dout <= 16'b0111001101100001;
        8'b01010010: dout <= 16'b0010110101110100;
        8'b01010011: dout <= 16'b0110000101111101;
        8'b01010100: dout <= 16'b0010100100100000;
        8'b01010110: dout <= 16'b0010000000100000;
        8'b01010111: dout <= 16'b0011000101110100;
        8'b01011000: dout <= 16'b0010111101100101;
        8'b01011001: dout <= 16'b0010100001011110;
        8'b01011010: dout <= 16'b0111001101111011;
        8'b01011011: dout <= 16'b0010110101100001;
        8'b01011100: dout <= 16'b0110000101110100;
        8'b01011101: dout <= 16'b0010100101111101;
        8'b01011110: dout <= 16'b0101111000100000;
        8'b01011111: dout <= 16'b0011001000100000;
        8'b01100001: dout <= 16'b0010000000100000;
        8'b01100010: dout <= 16'b0011000101011100;
        8'b01100011: dout <= 16'b0010111101100110;
        8'b01100100: dout <= 16'b0010100001110010;
        8'b01100101: dout <= 16'b0111001101100001;
        8'b01100110: dout <= 16'b0010110101100011;
        8'b01100111: dout <= 16'b0110000101111011;
        8'b01101000: dout <= 16'b0010100100110001;
        8'b01101001: dout <= 16'b0101111001111101;
        8'b01101010: dout <= 16'b0110111001111011;
        8'b01101011: dout <= 16'b0010000000101000;
        8'b01101100: dout <= 16'b0010000001101110;
        8'b01101101: dout <= 16'b0010000000101101;
        8'b01101110: dout <= 16'b0010000000110001;
        8'b01101111: dout <= 16'b0010000000101001;
        8'b01110000: dout <= 16'b0010000000100001;
        8'b01110001: dout <= 16'b0010000001111101;
        8'b01110010: dout <= 16'b0010000000100000;
        8'b01110011: dout <= 16'b0010000001110100;
        8'b01110100: dout <= 16'b0010000001011110;
        8'b01110101: dout <= 16'b0010000001111011;
        8'b01110110: dout <= 16'b0010000001101110;
        8'b01110111: dout <= 16'b0010000000101101;
        8'b01111000: dout <= 16'b0010000000110001;
        8'b01111001: dout <= 16'b0010000001111101;
        8'b01111010: dout <= 16'b0010000001100101;
        8'b01111011: dout <= 16'b0010000001011110;
        8'b01111100: dout <= 16'b0010000001111011;
        8'b01111101: dout <= 16'b0010000001100001;
        8'b01111110: dout <= 16'b0010000001110100;
        8'b01111111: dout <= 16'b0010000001111101;
        8'b10000001: dout <= 16'b0010000000100000;
        8'b10000010: dout <= 16'b0011000101011100;
        8'b10000011: dout <= 16'b0010111101100110;
        8'b10000100: dout <= 16'b0010100001110010;
        8'b10000101: dout <= 16'b0111001101100001;
        8'b10000110: dout <= 16'b0010110101100011;
        8'b10000111: dout <= 16'b0110000101111011;
        8'b10001000: dout <= 16'b0010100100110001;
        8'b10001001: dout <= 16'b0101111001111101;
        8'b10001010: dout <= 16'b0110101101111011;
        8'b10001011: dout <= 16'b0010000001011100;
        8'b10001100: dout <= 16'b0010000001000111;
        8'b10001101: dout <= 16'b0010000001100001;
        8'b10001110: dout <= 16'b0010000001101101;
        8'b10001111: dout <= 16'b0010000001101101;
        8'b10010000: dout <= 16'b0010000001100001;
        8'b10010001: dout <= 16'b0010000000101000;
        8'b10010010: dout <= 16'b0010000001101011;
        8'b10010011: dout <= 16'b0010000000101001;
        8'b10010100: dout <= 16'b0010000001111101;
        8'b10010101: dout <= 16'b0010000000100000;
        8'b10010110: dout <= 16'b0010000001110100;
        8'b10010111: dout <= 16'b0010000001011110;
        8'b10011000: dout <= 16'b0010000001111011;
        8'b10011001: dout <= 16'b0010000001101011;
        8'b10011010: dout <= 16'b0010000000101101;
        8'b10011011: dout <= 16'b0010000000110001;
        8'b10011100: dout <= 16'b0010000001111101;
        8'b10011101: dout <= 16'b0010000001100101;
        8'b10011110: dout <= 16'b0010000001011110;
        8'b10011111: dout <= 16'b0010000001111011;
        8'b10100000: dout <= 16'b0010000001100001;
        8'b10100001: dout <= 16'b0010000001110100;
        8'b10100010: dout <= 16'b0010000001111101;
        8'b10100100: dout <= 16'b0010000000100000;
        default: dout <= 16'b0010000000100000;
    endcase;
end

endmodule



module line_mapper(
//input wire clk,
//input wire rst,
input wire [7:0] line, 
output reg [15:0] addr);

//always @(posedge clk, posedge rst) begin
always @(line) begin
    // if (rst)
    //     addr <= 16'b0000001100000000;
    case(line)
    8'b00000000: addr <= 16'b0000001100000000;
    8'b00000001: addr <= 16'b0000010100000101;
    8'b00000010: addr <= 16'b0000111000001100;
    8'b00000011: addr <= 16'b0000111000011100;
    8'b00000100: addr <= 16'b0000110100101100;
    8'b00000101: addr <= 16'b0001000100111011;
    8'b00000110: addr <= 16'b0000011101001110;
    8'b00000111: addr <= 16'b0000100101010111;
    8'b00001000: addr <= 16'b0001111001100010;
    8'b00001001: addr <= 16'b0010000110000010;
    default: addr <= 16'b0000001100000000;
    endcase;
end

endmodule



